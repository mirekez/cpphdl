package MemWBint_int_0_0_State_pkg;

typedef struct packed {
    logic[8-1:0] _align0;
} MemWBint_int_0_0_State;


endpackage
