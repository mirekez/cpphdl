`default_nettype none

import Predef_pkg::*;
import DecodeFetchint_int_0_0_State_pkg::*;
import ExecuteCalcint_int_0_0_State_pkg::*;
import MakeBigStateDecodeFetchint_int_0_0_State_pkg::*;
import MemWBint_int_0_0_State_pkg::*;


module MemWBMemWBint_int_0_0_State_MakeBigStateDecodeFetchint_int_0_0_State_ExecuteCalcint_int_0_0_State_MemWBint_int_0_0_State #(
    parameter ID
,   parameter LENGTH
 )
 (
    input wire clk
,   input wire reset
,   input logic[31:0] mem_data_in
,   output logic[31:0] regs_data_out
,   output logic[7:0] regs_wr_id_out
,   output wire regs_write_out
,   input MakeBigStateDecodeFetchint_int_0_0_State[3-1:0] state_in
,   output MemWBint_int_0_0_State[1-1:0] state_out
);

    logic[31:0] regs_out_comb;
    logic regs_write_comb;
    MemWBint_int_0_0_State[1-1:0] state_reg;
    logic[63:0] i;

    task work (input logic reset);
    begin: work
        if (reset) begin
        end
    end
    endtask


    always @(posedge clk) begin
        work(reset);
    end

endmodule
