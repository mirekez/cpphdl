package Wb_pkg;

enum {
    WNONE,
    ALU,
    MEM,
    PC2,
    PC4
} Wb;


endpackage
