package ExecuteCalcint_int_0_0_State_pkg;

typedef struct packed {
    logic debug_branch_taken;
    logic[31:0] debug_branch_target;
    logic[31:0] debug_alu_b;
    logic[31:0] debug_alu_a;
    logic[31:0] alu_result;
} ExecuteCalcint_int_0_0_State;


endpackage
