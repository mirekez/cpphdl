package Mem_pkg;

enum {
    MNONE,
    LOAD,
    STORE
} Mem;


endpackage
