package Br_pkg;

enum {
    BNONE,
    BEQ,
    BNE,
    BLT,
    BGE,
    BLTU,
    BGEU,
    JAL,
    JALR,
    JR,
    BEQZ,
    BNEZ
} Br;


endpackage
