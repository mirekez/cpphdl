package MemWBint_int_0_0_State_pkg;

typedef struct packed {
    integer placeholder;
} MemWBint_int_0_0_State;


endpackage
