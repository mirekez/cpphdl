package Predef_pkg;

endpackage
