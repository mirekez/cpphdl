package MemWBint_int_0_0_State_pkg;

typedef struct packed {
    int dummy;
} MemWBint_int_0_0_State;


endpackage
