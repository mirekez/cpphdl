package Predef_pkg;

    parameter g_debug_en = 1;

endpackage
