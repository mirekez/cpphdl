package Alu_pkg;

enum {
    ANONE,
    ADD,
    SUB,
    AND,
    OR,
    XOR,
    SLL,
    SRL,
    SRA,
    SLT,
    SLTU,
    PASS,
    MUL,
    MULH,
    DIV,
    REM
} Alu;


endpackage
